module tb_integrated_designs ();

 //input signals
 reg tb_clk, tb_nrst;
 wire [3:0] tb_design_select;
 wire [33:0] tb_gpio_in, tb_gpio_oeb, tb_gpio_out;

 
    
endmodule