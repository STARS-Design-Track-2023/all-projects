VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO stopwatch
  CLASS BLOCK ;
  FOREIGN stopwatch ;
  ORIGIN 0.000 0.000 ;
  SIZE 154.895 BY 165.615 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 25.955 10.640 27.555 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 61.830 10.640 63.430 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 97.705 10.640 99.305 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 133.580 10.640 135.180 152.560 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 31.060 149.280 32.660 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 66.420 149.280 68.020 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 101.780 149.280 103.380 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 137.140 149.280 138.740 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 22.655 10.640 24.255 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 58.530 10.640 60.130 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 94.405 10.640 96.005 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 130.280 10.640 131.880 152.560 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 27.760 149.280 29.360 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 63.120 149.280 64.720 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 98.480 149.280 100.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 133.840 149.280 135.440 ;
    END
  END VPWR
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 37.440 4.000 38.040 ;
    END
  END clk
  PIN nrst
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 144.990 161.615 145.270 165.615 ;
    END
  END nrst
  PIN out_0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 74.150 0.000 74.430 4.000 ;
    END
  END out_0[0]
  PIN out_0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 48.390 161.615 48.670 165.615 ;
    END
  END out_0[1]
  PIN out_0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.840 4.000 58.440 ;
    END
  END out_0[2]
  PIN out_0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 150.895 54.440 154.895 55.040 ;
    END
  END out_0[3]
  PIN out_0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 87.030 161.615 87.310 165.615 ;
    END
  END out_0[4]
  PIN out_0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 151.430 0.000 151.710 4.000 ;
    END
  END out_0[5]
  PIN out_0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 150.895 95.240 154.895 95.840 ;
    END
  END out_0[6]
  PIN out_1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 132.110 0.000 132.390 4.000 ;
    END
  END out_1[0]
  PIN out_1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 150.895 115.640 154.895 116.240 ;
    END
  END out_1[1]
  PIN out_1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.040 4.000 17.640 ;
    END
  END out_1[2]
  PIN out_1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END out_1[3]
  PIN out_1[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 106.350 161.615 106.630 165.615 ;
    END
  END out_1[4]
  PIN out_1[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 125.670 161.615 125.950 165.615 ;
    END
  END out_1[5]
  PIN out_1[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.040 4.000 119.640 ;
    END
  END out_1[6]
  PIN out_2[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 29.070 161.615 29.350 165.615 ;
    END
  END out_2[0]
  PIN out_2[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 112.790 0.000 113.070 4.000 ;
    END
  END out_2[1]
  PIN out_2[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 139.440 4.000 140.040 ;
    END
  END out_2[2]
  PIN out_2[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 150.895 13.640 154.895 14.240 ;
    END
  END out_2[3]
  PIN out_2[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 16.190 0.000 16.470 4.000 ;
    END
  END out_2[4]
  PIN out_2[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 35.510 0.000 35.790 4.000 ;
    END
  END out_2[5]
  PIN out_2[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 9.750 161.615 10.030 165.615 ;
    END
  END out_2[6]
  PIN out_3[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 150.895 34.040 154.895 34.640 ;
    END
  END out_3[0]
  PIN out_3[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 54.830 0.000 55.110 4.000 ;
    END
  END out_3[1]
  PIN out_3[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 150.895 136.040 154.895 136.640 ;
    END
  END out_3[2]
  PIN out_3[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 150.895 156.440 154.895 157.040 ;
    END
  END out_3[3]
  PIN out_3[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 98.640 4.000 99.240 ;
    END
  END out_3[4]
  PIN out_3[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 67.710 161.615 67.990 165.615 ;
    END
  END out_3[5]
  PIN out_3[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 93.470 0.000 93.750 4.000 ;
    END
  END out_3[6]
  PIN pb_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.240 4.000 78.840 ;
    END
  END pb_0
  PIN pb_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 159.840 4.000 160.440 ;
    END
  END pb_1
  PIN time_done
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 150.895 74.840 154.895 75.440 ;
    END
  END time_done
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 149.040 152.405 ;
      LAYER met1 ;
        RECT 0.070 10.640 151.730 152.560 ;
      LAYER met2 ;
        RECT 0.100 161.335 9.470 162.250 ;
        RECT 10.310 161.335 28.790 162.250 ;
        RECT 29.630 161.335 48.110 162.250 ;
        RECT 48.950 161.335 67.430 162.250 ;
        RECT 68.270 161.335 86.750 162.250 ;
        RECT 87.590 161.335 106.070 162.250 ;
        RECT 106.910 161.335 125.390 162.250 ;
        RECT 126.230 161.335 144.710 162.250 ;
        RECT 145.550 161.335 151.700 162.250 ;
        RECT 0.100 4.280 151.700 161.335 ;
        RECT 0.650 4.000 15.910 4.280 ;
        RECT 16.750 4.000 35.230 4.280 ;
        RECT 36.070 4.000 54.550 4.280 ;
        RECT 55.390 4.000 73.870 4.280 ;
        RECT 74.710 4.000 93.190 4.280 ;
        RECT 94.030 4.000 112.510 4.280 ;
        RECT 113.350 4.000 131.830 4.280 ;
        RECT 132.670 4.000 151.150 4.280 ;
      LAYER met3 ;
        RECT 4.400 159.440 150.895 160.290 ;
        RECT 3.990 157.440 150.895 159.440 ;
        RECT 3.990 156.040 150.495 157.440 ;
        RECT 3.990 140.440 150.895 156.040 ;
        RECT 4.400 139.040 150.895 140.440 ;
        RECT 3.990 137.040 150.895 139.040 ;
        RECT 3.990 135.640 150.495 137.040 ;
        RECT 3.990 120.040 150.895 135.640 ;
        RECT 4.400 118.640 150.895 120.040 ;
        RECT 3.990 116.640 150.895 118.640 ;
        RECT 3.990 115.240 150.495 116.640 ;
        RECT 3.990 99.640 150.895 115.240 ;
        RECT 4.400 98.240 150.895 99.640 ;
        RECT 3.990 96.240 150.895 98.240 ;
        RECT 3.990 94.840 150.495 96.240 ;
        RECT 3.990 79.240 150.895 94.840 ;
        RECT 4.400 77.840 150.895 79.240 ;
        RECT 3.990 75.840 150.895 77.840 ;
        RECT 3.990 74.440 150.495 75.840 ;
        RECT 3.990 58.840 150.895 74.440 ;
        RECT 4.400 57.440 150.895 58.840 ;
        RECT 3.990 55.440 150.895 57.440 ;
        RECT 3.990 54.040 150.495 55.440 ;
        RECT 3.990 38.440 150.895 54.040 ;
        RECT 4.400 37.040 150.895 38.440 ;
        RECT 3.990 35.040 150.895 37.040 ;
        RECT 3.990 33.640 150.495 35.040 ;
        RECT 3.990 18.040 150.895 33.640 ;
        RECT 4.400 16.640 150.895 18.040 ;
        RECT 3.990 14.640 150.895 16.640 ;
        RECT 3.990 13.240 150.495 14.640 ;
        RECT 3.990 10.715 150.895 13.240 ;
      LAYER met4 ;
        RECT 73.895 60.015 94.005 117.465 ;
        RECT 96.405 60.015 97.305 117.465 ;
        RECT 99.705 60.015 99.985 117.465 ;
  END
END stopwatch
END LIBRARY

