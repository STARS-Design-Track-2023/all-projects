VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO silly_synthesizer
  CLASS BLOCK ;
  FOREIGN silly_synthesizer ;
  ORIGIN 0.000 0.000 ;
  SIZE 230.910 BY 241.630 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 24.340 10.640 25.940 228.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 177.940 10.640 179.540 228.720 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 30.030 225.180 31.630 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 183.210 225.180 184.810 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 228.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 228.720 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 26.730 225.180 28.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 179.910 225.180 181.510 ;
    END
  END VPWR
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 173.970 0.000 174.250 4.000 ;
    END
  END clk
  PIN cs
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 226.910 217.640 230.910 218.240 ;
    END
  END cs
  PIN gpio[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 209.390 237.630 209.670 241.630 ;
    END
  END gpio[0]
  PIN gpio[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 119.230 237.630 119.510 241.630 ;
    END
  END gpio[10]
  PIN gpio[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.240 4.000 44.840 ;
    END
  END gpio[11]
  PIN gpio[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 91.840 4.000 92.440 ;
    END
  END gpio[12]
  PIN gpio[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 226.910 30.640 230.910 31.240 ;
    END
  END gpio[13]
  PIN gpio[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 183.640 4.000 184.240 ;
    END
  END gpio[14]
  PIN gpio[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 226.910 170.040 230.910 170.640 ;
    END
  END gpio[15]
  PIN gpio[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END gpio[16]
  PIN gpio[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 41.950 0.000 42.230 4.000 ;
    END
  END gpio[1]
  PIN gpio[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 219.050 0.000 219.330 4.000 ;
    END
  END gpio[2]
  PIN gpio[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 87.030 0.000 87.310 4.000 ;
    END
  END gpio[3]
  PIN gpio[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 77.370 237.630 77.650 241.630 ;
    END
  END gpio[4]
  PIN gpio[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 226.910 122.440 230.910 123.040 ;
    END
  END gpio[5]
  PIN gpio[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 231.240 4.000 231.840 ;
    END
  END gpio[6]
  PIN gpio[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 164.310 237.630 164.590 241.630 ;
    END
  END gpio[7]
  PIN gpio[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 128.890 0.000 129.170 4.000 ;
    END
  END gpio[8]
  PIN gpio[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 136.040 4.000 136.640 ;
    END
  END gpio[9]
  PIN nrst
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 32.290 237.630 32.570 241.630 ;
    END
  END nrst
  PIN pwm
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 226.910 78.240 230.910 78.840 ;
    END
  END pwm
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 224.940 228.565 ;
      LAYER met1 ;
        RECT 0.070 10.640 225.790 228.720 ;
      LAYER met2 ;
        RECT 0.100 237.350 32.010 238.410 ;
        RECT 32.850 237.350 77.090 238.410 ;
        RECT 77.930 237.350 118.950 238.410 ;
        RECT 119.790 237.350 164.030 238.410 ;
        RECT 164.870 237.350 209.110 238.410 ;
        RECT 209.950 237.350 225.770 238.410 ;
        RECT 0.100 4.280 225.770 237.350 ;
        RECT 0.650 4.000 41.670 4.280 ;
        RECT 42.510 4.000 86.750 4.280 ;
        RECT 87.590 4.000 128.610 4.280 ;
        RECT 129.450 4.000 173.690 4.280 ;
        RECT 174.530 4.000 218.770 4.280 ;
        RECT 219.610 4.000 225.770 4.280 ;
      LAYER met3 ;
        RECT 4.400 230.840 226.910 231.690 ;
        RECT 4.000 218.640 226.910 230.840 ;
        RECT 4.000 217.240 226.510 218.640 ;
        RECT 4.000 184.640 226.910 217.240 ;
        RECT 4.400 183.240 226.910 184.640 ;
        RECT 4.000 171.040 226.910 183.240 ;
        RECT 4.000 169.640 226.510 171.040 ;
        RECT 4.000 137.040 226.910 169.640 ;
        RECT 4.400 135.640 226.910 137.040 ;
        RECT 4.000 123.440 226.910 135.640 ;
        RECT 4.000 122.040 226.510 123.440 ;
        RECT 4.000 92.840 226.910 122.040 ;
        RECT 4.400 91.440 226.910 92.840 ;
        RECT 4.000 79.240 226.910 91.440 ;
        RECT 4.000 77.840 226.510 79.240 ;
        RECT 4.000 45.240 226.910 77.840 ;
        RECT 4.400 43.840 226.910 45.240 ;
        RECT 4.000 31.640 226.910 43.840 ;
        RECT 4.000 30.240 226.510 31.640 ;
        RECT 4.000 10.715 226.910 30.240 ;
      LAYER met4 ;
        RECT 27.895 47.775 110.105 124.265 ;
  END
END silly_synthesizer
END LIBRARY

