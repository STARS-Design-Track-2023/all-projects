VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO Eighty_Twos
  CLASS BLOCK ;
  FOREIGN Eighty_Twos ;
  ORIGIN 0.000 0.000 ;
  SIZE 198.335 BY 209.055 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 24.340 10.640 25.940 196.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 177.940 10.640 179.540 196.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 30.030 192.980 31.630 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 183.210 192.980 184.810 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 196.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 196.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 26.730 192.980 28.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 179.910 192.980 181.510 ;
    END
  END VPWR
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 12.970 205.055 13.250 209.055 ;
    END
  END clk
  PIN cs
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 154.650 0.000 154.930 4.000 ;
    END
  END cs
  PIN gpi[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 176.840 4.000 177.440 ;
    END
  END gpi[0]
  PIN gpi[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 163.240 4.000 163.840 ;
    END
  END gpi[10]
  PIN gpi[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 194.335 119.040 198.335 119.640 ;
    END
  END gpi[11]
  PIN gpi[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.590 205.055 80.870 209.055 ;
    END
  END gpi[12]
  PIN gpi[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.290 205.055 193.570 209.055 ;
    END
  END gpi[13]
  PIN gpi[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 194.335 142.840 198.335 143.440 ;
    END
  END gpi[14]
  PIN gpi[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 194.335 37.440 198.335 38.040 ;
    END
  END gpi[15]
  PIN gpi[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 194.335 132.640 198.335 133.240 ;
    END
  END gpi[16]
  PIN gpi[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.990 0.000 145.270 4.000 ;
    END
  END gpi[17]
  PIN gpi[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 194.335 47.640 198.335 48.240 ;
    END
  END gpi[18]
  PIN gpi[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.040 4.000 34.640 ;
    END
  END gpi[19]
  PIN gpi[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 190.070 0.000 190.350 4.000 ;
    END
  END gpi[1]
  PIN gpi[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 194.335 23.840 198.335 24.440 ;
    END
  END gpi[20]
  PIN gpi[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.050 205.055 58.330 209.055 ;
    END
  END gpi[21]
  PIN gpi[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.030 0.000 87.310 4.000 ;
    END
  END gpi[22]
  PIN gpi[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 64.490 0.000 64.770 4.000 ;
    END
  END gpi[23]
  PIN gpi[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 153.040 4.000 153.640 ;
    END
  END gpi[24]
  PIN gpi[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.240 4.000 44.840 ;
    END
  END gpi[25]
  PIN gpi[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 194.335 156.440 198.335 157.040 ;
    END
  END gpi[26]
  PIN gpi[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 115.640 4.000 116.240 ;
    END
  END gpi[27]
  PIN gpi[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.570 0.000 109.850 4.000 ;
    END
  END gpi[28]
  PIN gpi[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 139.440 4.000 140.040 ;
    END
  END gpi[29]
  PIN gpi[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 194.335 166.640 198.335 167.240 ;
    END
  END gpi[2]
  PIN gpi[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 194.335 85.040 198.335 85.640 ;
    END
  END gpi[30]
  PIN gpi[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.210 205.055 148.490 209.055 ;
    END
  END gpi[31]
  PIN gpi[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.510 205.055 35.790 209.055 ;
    END
  END gpi[32]
  PIN gpi[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.950 0.000 42.230 4.000 ;
    END
  END gpi[33]
  PIN gpi[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 91.840 4.000 92.440 ;
    END
  END gpi[3]
  PIN gpi[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 20.440 4.000 21.040 ;
    END
  END gpi[4]
  PIN gpi[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 177.190 0.000 177.470 4.000 ;
    END
  END gpi[5]
  PIN gpi[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 103.130 205.055 103.410 209.055 ;
    END
  END gpi[6]
  PIN gpi[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 194.335 204.040 198.335 204.640 ;
    END
  END gpi[7]
  PIN gpi[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.530 0.000 167.810 4.000 ;
    END
  END gpi[8]
  PIN gpi[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.250 205.055 90.530 209.055 ;
    END
  END gpi[9]
  PIN gpo[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 194.335 13.640 198.335 14.240 ;
    END
  END gpo[0]
  PIN gpo[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 194.335 61.240 198.335 61.840 ;
    END
  END gpo[10]
  PIN gpo[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 122.450 0.000 122.730 4.000 ;
    END
  END gpo[11]
  PIN gpo[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 194.335 71.440 198.335 72.040 ;
    END
  END gpo[12]
  PIN gpo[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 125.670 205.055 125.950 209.055 ;
    END
  END gpo[13]
  PIN gpo[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 135.330 205.055 135.610 209.055 ;
    END
  END gpo[14]
  PIN gpo[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 0.090 205.055 0.370 209.055 ;
    END
  END gpo[15]
  PIN gpo[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END gpo[16]
  PIN gpo[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.240 4.000 129.840 ;
    END
  END gpo[17]
  PIN gpo[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 112.790 205.055 113.070 209.055 ;
    END
  END gpo[18]
  PIN gpo[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 157.870 205.055 158.150 209.055 ;
    END
  END gpo[19]
  PIN gpo[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 194.335 190.440 198.335 191.040 ;
    END
  END gpo[1]
  PIN gpo[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 67.710 205.055 67.990 209.055 ;
    END
  END gpo[20]
  PIN gpo[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 19.410 0.000 19.690 4.000 ;
    END
  END gpo[21]
  PIN gpo[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 9.750 0.000 10.030 4.000 ;
    END
  END gpo[22]
  PIN gpo[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 200.640 4.000 201.240 ;
    END
  END gpo[23]
  PIN gpo[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 180.410 205.055 180.690 209.055 ;
    END
  END gpo[24]
  PIN gpo[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 77.370 0.000 77.650 4.000 ;
    END
  END gpo[25]
  PIN gpo[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 194.335 180.240 198.335 180.840 ;
    END
  END gpo[26]
  PIN gpo[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 194.335 0.040 198.335 0.640 ;
    END
  END gpo[27]
  PIN gpo[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.840 4.000 58.440 ;
    END
  END gpo[28]
  PIN gpo[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.240 4.000 10.840 ;
    END
  END gpo[29]
  PIN gpo[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 32.290 0.000 32.570 4.000 ;
    END
  END gpo[2]
  PIN gpo[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 54.830 0.000 55.110 4.000 ;
    END
  END gpo[30]
  PIN gpo[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 105.440 4.000 106.040 ;
    END
  END gpo[31]
  PIN gpo[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 194.335 108.840 198.335 109.440 ;
    END
  END gpo[32]
  PIN gpo[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 99.910 0.000 100.190 4.000 ;
    END
  END gpo[33]
  PIN gpo[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 81.640 4.000 82.240 ;
    END
  END gpo[3]
  PIN gpo[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 170.750 205.055 171.030 209.055 ;
    END
  END gpo[4]
  PIN gpo[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 22.630 205.055 22.910 209.055 ;
    END
  END gpo[5]
  PIN gpo[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 45.170 205.055 45.450 209.055 ;
    END
  END gpo[6]
  PIN gpo[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 132.110 0.000 132.390 4.000 ;
    END
  END gpo[7]
  PIN gpo[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.040 4.000 68.640 ;
    END
  END gpo[8]
  PIN gpo[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 187.040 4.000 187.640 ;
    END
  END gpo[9]
  PIN nrst
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 194.335 95.240 198.335 95.840 ;
    END
  END nrst
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 192.740 195.925 ;
      LAYER met1 ;
        RECT 0.070 10.640 192.740 196.080 ;
      LAYER met2 ;
        RECT 0.650 204.775 12.690 205.770 ;
        RECT 13.530 204.775 22.350 205.770 ;
        RECT 23.190 204.775 35.230 205.770 ;
        RECT 36.070 204.775 44.890 205.770 ;
        RECT 45.730 204.775 57.770 205.770 ;
        RECT 58.610 204.775 67.430 205.770 ;
        RECT 68.270 204.775 80.310 205.770 ;
        RECT 81.150 204.775 89.970 205.770 ;
        RECT 90.810 204.775 102.850 205.770 ;
        RECT 103.690 204.775 112.510 205.770 ;
        RECT 113.350 204.775 125.390 205.770 ;
        RECT 126.230 204.775 135.050 205.770 ;
        RECT 135.890 204.775 147.930 205.770 ;
        RECT 148.770 204.775 157.590 205.770 ;
        RECT 158.430 204.775 170.470 205.770 ;
        RECT 171.310 204.775 180.130 205.770 ;
        RECT 180.970 204.775 192.650 205.770 ;
        RECT 0.100 4.280 192.650 204.775 ;
        RECT 0.650 0.155 9.470 4.280 ;
        RECT 10.310 0.155 19.130 4.280 ;
        RECT 19.970 0.155 32.010 4.280 ;
        RECT 32.850 0.155 41.670 4.280 ;
        RECT 42.510 0.155 54.550 4.280 ;
        RECT 55.390 0.155 64.210 4.280 ;
        RECT 65.050 0.155 77.090 4.280 ;
        RECT 77.930 0.155 86.750 4.280 ;
        RECT 87.590 0.155 99.630 4.280 ;
        RECT 100.470 0.155 109.290 4.280 ;
        RECT 110.130 0.155 122.170 4.280 ;
        RECT 123.010 0.155 131.830 4.280 ;
        RECT 132.670 0.155 144.710 4.280 ;
        RECT 145.550 0.155 154.370 4.280 ;
        RECT 155.210 0.155 167.250 4.280 ;
        RECT 168.090 0.155 176.910 4.280 ;
        RECT 177.750 0.155 189.790 4.280 ;
        RECT 190.630 0.155 192.650 4.280 ;
      LAYER met3 ;
        RECT 4.000 203.640 193.935 204.505 ;
        RECT 4.000 201.640 194.335 203.640 ;
        RECT 4.400 200.240 194.335 201.640 ;
        RECT 4.000 191.440 194.335 200.240 ;
        RECT 4.000 190.040 193.935 191.440 ;
        RECT 4.000 188.040 194.335 190.040 ;
        RECT 4.400 186.640 194.335 188.040 ;
        RECT 4.000 181.240 194.335 186.640 ;
        RECT 4.000 179.840 193.935 181.240 ;
        RECT 4.000 177.840 194.335 179.840 ;
        RECT 4.400 176.440 194.335 177.840 ;
        RECT 4.000 167.640 194.335 176.440 ;
        RECT 4.000 166.240 193.935 167.640 ;
        RECT 4.000 164.240 194.335 166.240 ;
        RECT 4.400 162.840 194.335 164.240 ;
        RECT 4.000 157.440 194.335 162.840 ;
        RECT 4.000 156.040 193.935 157.440 ;
        RECT 4.000 154.040 194.335 156.040 ;
        RECT 4.400 152.640 194.335 154.040 ;
        RECT 4.000 143.840 194.335 152.640 ;
        RECT 4.000 142.440 193.935 143.840 ;
        RECT 4.000 140.440 194.335 142.440 ;
        RECT 4.400 139.040 194.335 140.440 ;
        RECT 4.000 133.640 194.335 139.040 ;
        RECT 4.000 132.240 193.935 133.640 ;
        RECT 4.000 130.240 194.335 132.240 ;
        RECT 4.400 128.840 194.335 130.240 ;
        RECT 4.000 120.040 194.335 128.840 ;
        RECT 4.000 118.640 193.935 120.040 ;
        RECT 4.000 116.640 194.335 118.640 ;
        RECT 4.400 115.240 194.335 116.640 ;
        RECT 4.000 109.840 194.335 115.240 ;
        RECT 4.000 108.440 193.935 109.840 ;
        RECT 4.000 106.440 194.335 108.440 ;
        RECT 4.400 105.040 194.335 106.440 ;
        RECT 4.000 96.240 194.335 105.040 ;
        RECT 4.000 94.840 193.935 96.240 ;
        RECT 4.000 92.840 194.335 94.840 ;
        RECT 4.400 91.440 194.335 92.840 ;
        RECT 4.000 86.040 194.335 91.440 ;
        RECT 4.000 84.640 193.935 86.040 ;
        RECT 4.000 82.640 194.335 84.640 ;
        RECT 4.400 81.240 194.335 82.640 ;
        RECT 4.000 72.440 194.335 81.240 ;
        RECT 4.000 71.040 193.935 72.440 ;
        RECT 4.000 69.040 194.335 71.040 ;
        RECT 4.400 67.640 194.335 69.040 ;
        RECT 4.000 62.240 194.335 67.640 ;
        RECT 4.000 60.840 193.935 62.240 ;
        RECT 4.000 58.840 194.335 60.840 ;
        RECT 4.400 57.440 194.335 58.840 ;
        RECT 4.000 48.640 194.335 57.440 ;
        RECT 4.000 47.240 193.935 48.640 ;
        RECT 4.000 45.240 194.335 47.240 ;
        RECT 4.400 43.840 194.335 45.240 ;
        RECT 4.000 38.440 194.335 43.840 ;
        RECT 4.000 37.040 193.935 38.440 ;
        RECT 4.000 35.040 194.335 37.040 ;
        RECT 4.400 33.640 194.335 35.040 ;
        RECT 4.000 24.840 194.335 33.640 ;
        RECT 4.000 23.440 193.935 24.840 ;
        RECT 4.000 21.440 194.335 23.440 ;
        RECT 4.400 20.040 194.335 21.440 ;
        RECT 4.000 14.640 194.335 20.040 ;
        RECT 4.000 13.240 193.935 14.640 ;
        RECT 4.000 11.240 194.335 13.240 ;
        RECT 4.400 9.840 194.335 11.240 ;
        RECT 4.000 1.040 194.335 9.840 ;
        RECT 4.000 0.175 193.935 1.040 ;
      LAYER met4 ;
        RECT 49.055 13.095 174.240 194.305 ;
        RECT 176.640 13.095 177.540 194.305 ;
        RECT 179.940 13.095 180.945 194.305 ;
  END
END Eighty_Twos
END LIBRARY

