VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO Synthia
  CLASS BLOCK ;
  FOREIGN Synthia ;
  ORIGIN 0.000 0.000 ;
  SIZE 266.535 BY 277.255 ;
  PIN PWM_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 262.535 27.240 266.535 27.840 ;
    END
  END PWM_o
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 24.340 10.640 25.940 264.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 177.940 10.640 179.540 264.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 30.030 261.060 31.630 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 183.210 261.060 184.810 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 264.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 264.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 26.730 261.060 28.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 179.910 261.060 181.510 ;
    END
  END VPWR
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 262.535 214.240 266.535 214.840 ;
    END
  END clk
  PIN modes
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 148.210 273.255 148.490 277.255 ;
    END
  END modes
  PIN octaves
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 177.190 0.000 177.470 4.000 ;
    END
  END octaves
  PIN pb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 248.240 4.000 248.840 ;
    END
  END pb[0]
  PIN pb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 87.030 273.255 87.310 277.255 ;
    END
  END pb[10]
  PIN pb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END pb[11]
  PIN pb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 264.130 273.255 264.410 277.255 ;
    END
  END pb[12]
  PIN pb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 235.150 0.000 235.430 4.000 ;
    END
  END pb[1]
  PIN pb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 58.050 0.000 58.330 4.000 ;
    END
  END pb[2]
  PIN pb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.240 4.000 61.840 ;
    END
  END pb[3]
  PIN pb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 262.535 153.040 266.535 153.640 ;
    END
  END pb[4]
  PIN pb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 122.440 4.000 123.040 ;
    END
  END pb[5]
  PIN pb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 206.170 273.255 206.450 277.255 ;
    END
  END pb[6]
  PIN pb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 116.010 0.000 116.290 4.000 ;
    END
  END pb[7]
  PIN pb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 183.640 4.000 184.240 ;
    END
  END pb[8]
  PIN pb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 29.070 273.255 29.350 277.255 ;
    END
  END pb[9]
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 262.535 91.840 266.535 92.440 ;
    END
  END reset
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 260.820 263.925 ;
      LAYER met1 ;
        RECT 0.070 10.640 264.430 264.080 ;
      LAYER met2 ;
        RECT 0.100 272.975 28.790 273.255 ;
        RECT 29.630 272.975 86.750 273.255 ;
        RECT 87.590 272.975 147.930 273.255 ;
        RECT 148.770 272.975 205.890 273.255 ;
        RECT 206.730 272.975 263.850 273.255 ;
        RECT 0.100 4.280 264.400 272.975 ;
        RECT 0.650 4.000 57.770 4.280 ;
        RECT 58.610 4.000 115.730 4.280 ;
        RECT 116.570 4.000 176.910 4.280 ;
        RECT 177.750 4.000 234.870 4.280 ;
        RECT 235.710 4.000 264.400 4.280 ;
      LAYER met3 ;
        RECT 4.000 249.240 262.535 264.005 ;
        RECT 4.400 247.840 262.535 249.240 ;
        RECT 4.000 215.240 262.535 247.840 ;
        RECT 4.000 213.840 262.135 215.240 ;
        RECT 4.000 184.640 262.535 213.840 ;
        RECT 4.400 183.240 262.535 184.640 ;
        RECT 4.000 154.040 262.535 183.240 ;
        RECT 4.000 152.640 262.135 154.040 ;
        RECT 4.000 123.440 262.535 152.640 ;
        RECT 4.400 122.040 262.535 123.440 ;
        RECT 4.000 92.840 262.535 122.040 ;
        RECT 4.000 91.440 262.135 92.840 ;
        RECT 4.000 62.240 262.535 91.440 ;
        RECT 4.400 60.840 262.535 62.240 ;
        RECT 4.000 28.240 262.535 60.840 ;
        RECT 4.000 26.840 262.135 28.240 ;
        RECT 4.000 10.715 262.535 26.840 ;
      LAYER met4 ;
        RECT 66.535 12.415 174.240 241.225 ;
        RECT 176.640 12.415 177.540 241.225 ;
        RECT 179.940 12.415 211.305 241.225 ;
  END
END Synthia
END LIBRARY

