VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sass_synth
  CLASS BLOCK ;
  FOREIGN sass_synth ;
  ORIGIN 0.000 0.000 ;
  SIZE 366.095 BY 376.815 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 24.340 10.640 25.940 364.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 177.940 10.640 179.540 364.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 331.540 10.640 333.140 364.720 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 30.030 360.420 31.630 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 183.210 360.420 184.810 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 336.390 360.420 337.990 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 364.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 364.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 364.720 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 26.730 360.420 28.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 179.910 360.420 181.510 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 333.090 360.420 334.690 ;
    END
  END VPWR
  PIN beat_led[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 80.590 0.000 80.870 4.000 ;
    END
  END beat_led[0]
  PIN beat_led[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 227.840 4.000 228.440 ;
    END
  END beat_led[1]
  PIN beat_led[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 299.550 0.000 299.830 4.000 ;
    END
  END beat_led[2]
  PIN beat_led[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 22.630 372.815 22.910 376.815 ;
    END
  END beat_led[3]
  PIN beat_led[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 362.095 187.040 366.095 187.640 ;
    END
  END beat_led[4]
  PIN beat_led[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 270.570 0.000 270.850 4.000 ;
    END
  END beat_led[5]
  PIN beat_led[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 215.830 0.000 216.110 4.000 ;
    END
  END beat_led[6]
  PIN beat_led[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 285.640 4.000 286.240 ;
    END
  END beat_led[7]
  PIN cs
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 374.040 4.000 374.640 ;
    END
  END cs
  PIN hwclk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 362.095 44.240 366.095 44.840 ;
    END
  END hwclk
  PIN mode_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 241.590 372.815 241.870 376.815 ;
    END
  END mode_out[0]
  PIN mode_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 362.095 13.640 366.095 14.240 ;
    END
  END mode_out[1]
  PIN multi[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 296.330 372.815 296.610 376.815 ;
    END
  END multi[0]
  PIN multi[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 362.095 71.440 366.095 72.040 ;
    END
  END multi[1]
  PIN multi[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 51.610 372.815 51.890 376.815 ;
    END
  END multi[2]
  PIN multi[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 362.095 102.040 366.095 102.640 ;
    END
  END multi[3]
  PIN n_rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 258.440 4.000 259.040 ;
    END
  END n_rst
  PIN note1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 362.095 333.240 366.095 333.840 ;
    END
  END note1[0]
  PIN note1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.240 4.000 112.840 ;
    END
  END note1[1]
  PIN note1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 170.040 4.000 170.640 ;
    END
  END note1[2]
  PIN note1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 316.240 4.000 316.840 ;
    END
  END note1[3]
  PIN note2[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 354.290 0.000 354.570 4.000 ;
    END
  END note2[0]
  PIN note2[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 200.640 4.000 201.240 ;
    END
  END note2[1]
  PIN note2[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 362.095 275.440 366.095 276.040 ;
    END
  END note2[2]
  PIN note2[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.440 4.000 55.040 ;
    END
  END note2[3]
  PIN note3[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 215.830 372.815 216.110 376.815 ;
    END
  END note3[0]
  PIN note3[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.040 4.000 85.640 ;
    END
  END note3[1]
  PIN note3[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 362.095 360.440 366.095 361.040 ;
    END
  END note3[2]
  PIN note3[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 161.090 372.815 161.370 376.815 ;
    END
  END note3[3]
  PIN note4[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 362.095 217.640 366.095 218.240 ;
    END
  END note4[0]
  PIN note4[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 270.570 372.815 270.850 376.815 ;
    END
  END note4[1]
  PIN note4[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 25.850 0.000 26.130 4.000 ;
    END
  END note4[2]
  PIN note4[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END note4[3]
  PIN piano_keys[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 106.350 372.815 106.630 376.815 ;
    END
  END piano_keys[0]
  PIN piano_keys[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 362.095 302.640 366.095 303.240 ;
    END
  END piano_keys[10]
  PIN piano_keys[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 135.330 0.000 135.610 4.000 ;
    END
  END piano_keys[11]
  PIN piano_keys[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 362.095 244.840 366.095 245.440 ;
    END
  END piano_keys[12]
  PIN piano_keys[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 325.310 0.000 325.590 4.000 ;
    END
  END piano_keys[13]
  PIN piano_keys[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 186.850 372.815 187.130 376.815 ;
    END
  END piano_keys[14]
  PIN piano_keys[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 362.095 129.240 366.095 129.840 ;
    END
  END piano_keys[1]
  PIN piano_keys[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 51.610 0.000 51.890 4.000 ;
    END
  END piano_keys[2]
  PIN piano_keys[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 106.350 0.000 106.630 4.000 ;
    END
  END piano_keys[3]
  PIN piano_keys[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 161.090 0.000 161.370 4.000 ;
    END
  END piano_keys[4]
  PIN piano_keys[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.240 4.000 27.840 ;
    END
  END piano_keys[5]
  PIN piano_keys[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 190.070 0.000 190.350 4.000 ;
    END
  END piano_keys[6]
  PIN piano_keys[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 351.070 372.815 351.350 376.815 ;
    END
  END piano_keys[7]
  PIN piano_keys[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 325.310 372.815 325.590 376.815 ;
    END
  END piano_keys[8]
  PIN piano_keys[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 77.370 372.815 77.650 376.815 ;
    END
  END piano_keys[9]
  PIN pwm_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 132.110 372.815 132.390 376.815 ;
    END
  END pwm_o
  PIN seq_led_on
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 244.810 0.000 245.090 4.000 ;
    END
  END seq_led_on
  PIN seq_play
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 142.840 4.000 143.440 ;
    END
  END seq_play
  PIN seq_power
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 343.440 4.000 344.040 ;
    END
  END seq_power
  PIN tempo_select
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 362.095 159.840 366.095 160.440 ;
    END
  END tempo_select
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 360.180 364.565 ;
      LAYER met1 ;
        RECT 0.070 9.960 361.030 364.720 ;
      LAYER met2 ;
        RECT 0.100 372.535 22.350 374.525 ;
        RECT 23.190 372.535 51.330 374.525 ;
        RECT 52.170 372.535 77.090 374.525 ;
        RECT 77.930 372.535 106.070 374.525 ;
        RECT 106.910 372.535 131.830 374.525 ;
        RECT 132.670 372.535 160.810 374.525 ;
        RECT 161.650 372.535 186.570 374.525 ;
        RECT 187.410 372.535 215.550 374.525 ;
        RECT 216.390 372.535 241.310 374.525 ;
        RECT 242.150 372.535 270.290 374.525 ;
        RECT 271.130 372.535 296.050 374.525 ;
        RECT 296.890 372.535 325.030 374.525 ;
        RECT 325.870 372.535 350.790 374.525 ;
        RECT 351.630 372.535 361.010 374.525 ;
        RECT 0.100 4.280 361.010 372.535 ;
        RECT 0.650 3.670 25.570 4.280 ;
        RECT 26.410 3.670 51.330 4.280 ;
        RECT 52.170 3.670 80.310 4.280 ;
        RECT 81.150 3.670 106.070 4.280 ;
        RECT 106.910 3.670 135.050 4.280 ;
        RECT 135.890 3.670 160.810 4.280 ;
        RECT 161.650 3.670 189.790 4.280 ;
        RECT 190.630 3.670 215.550 4.280 ;
        RECT 216.390 3.670 244.530 4.280 ;
        RECT 245.370 3.670 270.290 4.280 ;
        RECT 271.130 3.670 299.270 4.280 ;
        RECT 300.110 3.670 325.030 4.280 ;
        RECT 325.870 3.670 354.010 4.280 ;
        RECT 354.850 3.670 361.010 4.280 ;
      LAYER met3 ;
        RECT 4.400 373.640 362.095 374.505 ;
        RECT 3.990 361.440 362.095 373.640 ;
        RECT 3.990 360.040 361.695 361.440 ;
        RECT 3.990 344.440 362.095 360.040 ;
        RECT 4.400 343.040 362.095 344.440 ;
        RECT 3.990 334.240 362.095 343.040 ;
        RECT 3.990 332.840 361.695 334.240 ;
        RECT 3.990 317.240 362.095 332.840 ;
        RECT 4.400 315.840 362.095 317.240 ;
        RECT 3.990 303.640 362.095 315.840 ;
        RECT 3.990 302.240 361.695 303.640 ;
        RECT 3.990 286.640 362.095 302.240 ;
        RECT 4.400 285.240 362.095 286.640 ;
        RECT 3.990 276.440 362.095 285.240 ;
        RECT 3.990 275.040 361.695 276.440 ;
        RECT 3.990 259.440 362.095 275.040 ;
        RECT 4.400 258.040 362.095 259.440 ;
        RECT 3.990 245.840 362.095 258.040 ;
        RECT 3.990 244.440 361.695 245.840 ;
        RECT 3.990 228.840 362.095 244.440 ;
        RECT 4.400 227.440 362.095 228.840 ;
        RECT 3.990 218.640 362.095 227.440 ;
        RECT 3.990 217.240 361.695 218.640 ;
        RECT 3.990 201.640 362.095 217.240 ;
        RECT 4.400 200.240 362.095 201.640 ;
        RECT 3.990 188.040 362.095 200.240 ;
        RECT 3.990 186.640 361.695 188.040 ;
        RECT 3.990 171.040 362.095 186.640 ;
        RECT 4.400 169.640 362.095 171.040 ;
        RECT 3.990 160.840 362.095 169.640 ;
        RECT 3.990 159.440 361.695 160.840 ;
        RECT 3.990 143.840 362.095 159.440 ;
        RECT 4.400 142.440 362.095 143.840 ;
        RECT 3.990 130.240 362.095 142.440 ;
        RECT 3.990 128.840 361.695 130.240 ;
        RECT 3.990 113.240 362.095 128.840 ;
        RECT 4.400 111.840 362.095 113.240 ;
        RECT 3.990 103.040 362.095 111.840 ;
        RECT 3.990 101.640 361.695 103.040 ;
        RECT 3.990 86.040 362.095 101.640 ;
        RECT 4.400 84.640 362.095 86.040 ;
        RECT 3.990 72.440 362.095 84.640 ;
        RECT 3.990 71.040 361.695 72.440 ;
        RECT 3.990 55.440 362.095 71.040 ;
        RECT 4.400 54.040 362.095 55.440 ;
        RECT 3.990 45.240 362.095 54.040 ;
        RECT 3.990 43.840 361.695 45.240 ;
        RECT 3.990 28.240 362.095 43.840 ;
        RECT 4.400 26.840 362.095 28.240 ;
        RECT 3.990 14.640 362.095 26.840 ;
        RECT 3.990 13.240 361.695 14.640 ;
        RECT 3.990 10.715 362.095 13.240 ;
      LAYER met4 ;
        RECT 95.975 58.655 174.240 363.625 ;
        RECT 176.640 58.655 177.540 363.625 ;
        RECT 179.940 58.655 327.840 363.625 ;
        RECT 330.240 58.655 331.140 363.625 ;
        RECT 333.540 58.655 348.385 363.625 ;
      LAYER met5 ;
        RECT 144.100 186.410 209.180 206.500 ;
        RECT 144.100 140.300 209.180 178.310 ;
  END
END sass_synth
END LIBRARY

