VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO top_asic
  CLASS BLOCK ;
  FOREIGN top_asic ;
  ORIGIN 0.000 0.000 ;
  SIZE 435.755 BY 446.475 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 24.340 10.640 25.940 435.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 177.940 10.640 179.540 435.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 331.540 10.640 333.140 435.440 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 30.030 430.340 31.630 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 183.210 430.340 184.810 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 336.390 430.340 337.990 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 435.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 435.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 435.440 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 26.730 430.340 28.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 179.910 430.340 181.510 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 333.090 430.340 334.690 ;
    END
  END VPWR
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 431.755 81.640 435.755 82.240 ;
    END
  END clk
  PIN mode_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 434.790 442.475 435.070 446.475 ;
    END
  END mode_out[0]
  PIN mode_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 264.130 442.475 264.410 446.475 ;
    END
  END mode_out[1]
  PIN pb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 170.750 0.000 171.030 4.000 ;
    END
  END pb[0]
  PIN pb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 431.755 357.040 435.755 357.640 ;
    END
  END pb[10]
  PIN pb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 431.570 0.000 431.850 4.000 ;
    END
  END pb[11]
  PIN pb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 363.840 4.000 364.440 ;
    END
  END pb[12]
  PIN pb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 177.190 442.475 177.470 446.475 ;
    END
  END pb[13]
  PIN pb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END pb[14]
  PIN pb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 90.250 442.475 90.530 446.475 ;
    END
  END pb[1]
  PIN pb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 344.630 0.000 344.910 4.000 ;
    END
  END pb[2]
  PIN pb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 83.810 0.000 84.090 4.000 ;
    END
  END pb[3]
  PIN pb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 88.440 4.000 89.040 ;
    END
  END pb[4]
  PIN pb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 431.755 265.240 435.755 265.840 ;
    END
  END pb[5]
  PIN pb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 180.240 4.000 180.840 ;
    END
  END pb[6]
  PIN pb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 351.070 442.475 351.350 446.475 ;
    END
  END pb[7]
  PIN pb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 257.690 0.000 257.970 4.000 ;
    END
  END pb[8]
  PIN pb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 272.040 4.000 272.640 ;
    END
  END pb[9]
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 3.310 442.475 3.590 446.475 ;
    END
  END reset
  PIN sigout
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 431.755 173.440 435.755 174.040 ;
    END
  END sigout
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 430.100 435.285 ;
      LAYER met1 ;
        RECT 0.070 10.640 435.090 435.440 ;
      LAYER met2 ;
        RECT 0.100 442.195 3.030 442.475 ;
        RECT 3.870 442.195 89.970 442.475 ;
        RECT 90.810 442.195 176.910 442.475 ;
        RECT 177.750 442.195 263.850 442.475 ;
        RECT 264.690 442.195 350.790 442.475 ;
        RECT 351.630 442.195 434.510 442.475 ;
        RECT 0.100 4.280 435.060 442.195 ;
        RECT 0.650 3.670 83.530 4.280 ;
        RECT 84.370 3.670 170.470 4.280 ;
        RECT 171.310 3.670 257.410 4.280 ;
        RECT 258.250 3.670 344.350 4.280 ;
        RECT 345.190 3.670 431.290 4.280 ;
        RECT 432.130 3.670 435.060 4.280 ;
      LAYER met3 ;
        RECT 3.990 364.840 431.755 435.365 ;
        RECT 4.400 363.440 431.755 364.840 ;
        RECT 3.990 358.040 431.755 363.440 ;
        RECT 3.990 356.640 431.355 358.040 ;
        RECT 3.990 273.040 431.755 356.640 ;
        RECT 4.400 271.640 431.755 273.040 ;
        RECT 3.990 266.240 431.755 271.640 ;
        RECT 3.990 264.840 431.355 266.240 ;
        RECT 3.990 181.240 431.755 264.840 ;
        RECT 4.400 179.840 431.755 181.240 ;
        RECT 3.990 174.440 431.755 179.840 ;
        RECT 3.990 173.040 431.355 174.440 ;
        RECT 3.990 89.440 431.755 173.040 ;
        RECT 4.400 88.040 431.755 89.440 ;
        RECT 3.990 82.640 431.755 88.040 ;
        RECT 3.990 81.240 431.355 82.640 ;
        RECT 3.990 10.715 431.755 81.240 ;
      LAYER met4 ;
        RECT 68.375 39.615 174.240 425.505 ;
        RECT 176.640 39.615 177.540 425.505 ;
        RECT 179.940 39.615 327.840 425.505 ;
        RECT 330.240 39.615 331.140 425.505 ;
        RECT 333.540 39.615 379.665 425.505 ;
      LAYER met5 ;
        RECT 136.740 186.410 374.780 308.500 ;
        RECT 136.740 147.100 374.780 178.310 ;
  END
END top_asic
END LIBRARY

