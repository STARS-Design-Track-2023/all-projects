VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO Guitar_Villains
  CLASS BLOCK ;
  FOREIGN Guitar_Villains ;
  ORIGIN 0.000 0.000 ;
  SIZE 315.970 BY 326.690 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 24.340 10.640 25.940 315.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 177.940 10.640 179.540 315.760 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 30.030 310.280 31.630 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 183.210 310.280 184.810 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 315.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 315.760 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 26.730 310.280 28.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 179.910 310.280 181.510 ;
    END
  END VPWR
  PIN bottom_row[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 167.530 0.000 167.810 4.000 ;
    END
  END bottom_row[0]
  PIN bottom_row[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 302.770 0.000 303.050 4.000 ;
    END
  END bottom_row[1]
  PIN bottom_row[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 61.270 322.690 61.550 326.690 ;
    END
  END bottom_row[2]
  PIN bottom_row[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 267.350 322.690 267.630 326.690 ;
    END
  END bottom_row[3]
  PIN bottom_row[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 105.440 4.000 106.040 ;
    END
  END bottom_row[4]
  PIN bottom_row[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 99.910 0.000 100.190 4.000 ;
    END
  END bottom_row[5]
  PIN bottom_row[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 270.570 0.000 270.850 4.000 ;
    END
  END bottom_row[6]
  PIN button[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 231.930 322.690 232.210 326.690 ;
    END
  END button[0]
  PIN button[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 214.240 4.000 214.840 ;
    END
  END button[1]
  PIN button[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 311.970 200.640 315.970 201.240 ;
    END
  END button[2]
  PIN button[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 199.730 322.690 200.010 326.690 ;
    END
  END button[3]
  PIN chip_select
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 285.640 4.000 286.240 ;
    END
  END chip_select
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 248.240 4.000 248.840 ;
    END
  END clk
  PIN green_disp
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 311.970 20.440 315.970 21.040 ;
    END
  END green_disp
  PIN n_rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 311.970 163.240 315.970 163.840 ;
    END
  END n_rst
  PIN red_disp
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 311.970 234.640 315.970 235.240 ;
    END
  END red_disp
  PIN ss0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END ss0[0]
  PIN ss0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 164.310 322.690 164.590 326.690 ;
    END
  END ss0[1]
  PIN ss0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.040 4.000 34.640 ;
    END
  END ss0[2]
  PIN ss0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 96.690 322.690 96.970 326.690 ;
    END
  END ss0[3]
  PIN ss0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 29.070 322.690 29.350 326.690 ;
    END
  END ss0[4]
  PIN ss0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 235.150 0.000 235.430 4.000 ;
    END
  END ss0[5]
  PIN ss0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 299.550 322.690 299.830 326.690 ;
    END
  END ss0[6]
  PIN ss1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 311.970 54.440 315.970 55.040 ;
    END
  END ss1[0]
  PIN ss1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 32.290 0.000 32.570 4.000 ;
    END
  END ss1[1]
  PIN ss1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 67.710 0.000 67.990 4.000 ;
    END
  END ss1[2]
  PIN ss1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 71.440 4.000 72.040 ;
    END
  END ss1[3]
  PIN ss1[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 311.970 91.840 315.970 92.440 ;
    END
  END ss1[4]
  PIN ss1[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 135.330 0.000 135.610 4.000 ;
    END
  END ss1[5]
  PIN ss1[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 311.970 272.040 315.970 272.640 ;
    END
  END ss1[6]
  PIN top_row[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 311.970 306.040 315.970 306.640 ;
    END
  END top_row[0]
  PIN top_row[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 176.840 4.000 177.440 ;
    END
  END top_row[1]
  PIN top_row[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 132.110 322.690 132.390 326.690 ;
    END
  END top_row[2]
  PIN top_row[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 202.950 0.000 203.230 4.000 ;
    END
  END top_row[3]
  PIN top_row[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 142.840 4.000 143.440 ;
    END
  END top_row[4]
  PIN top_row[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 319.640 4.000 320.240 ;
    END
  END top_row[5]
  PIN top_row[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 311.970 129.240 315.970 129.840 ;
    END
  END top_row[6]
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 310.040 315.605 ;
      LAYER met1 ;
        RECT 0.070 10.640 310.430 315.760 ;
      LAYER met2 ;
        RECT 0.100 322.410 28.790 323.410 ;
        RECT 29.630 322.410 60.990 323.410 ;
        RECT 61.830 322.410 96.410 323.410 ;
        RECT 97.250 322.410 131.830 323.410 ;
        RECT 132.670 322.410 164.030 323.410 ;
        RECT 164.870 322.410 199.450 323.410 ;
        RECT 200.290 322.410 231.650 323.410 ;
        RECT 232.490 322.410 267.070 323.410 ;
        RECT 267.910 322.410 299.270 323.410 ;
        RECT 300.110 322.410 310.410 323.410 ;
        RECT 0.100 4.280 310.410 322.410 ;
        RECT 0.650 3.670 32.010 4.280 ;
        RECT 32.850 3.670 67.430 4.280 ;
        RECT 68.270 3.670 99.630 4.280 ;
        RECT 100.470 3.670 135.050 4.280 ;
        RECT 135.890 3.670 167.250 4.280 ;
        RECT 168.090 3.670 202.670 4.280 ;
        RECT 203.510 3.670 234.870 4.280 ;
        RECT 235.710 3.670 270.290 4.280 ;
        RECT 271.130 3.670 302.490 4.280 ;
        RECT 303.330 3.670 310.410 4.280 ;
      LAYER met3 ;
        RECT 4.400 319.240 311.970 320.090 ;
        RECT 4.000 307.040 311.970 319.240 ;
        RECT 4.000 305.640 311.570 307.040 ;
        RECT 4.000 286.640 311.970 305.640 ;
        RECT 4.400 285.240 311.970 286.640 ;
        RECT 4.000 273.040 311.970 285.240 ;
        RECT 4.000 271.640 311.570 273.040 ;
        RECT 4.000 249.240 311.970 271.640 ;
        RECT 4.400 247.840 311.970 249.240 ;
        RECT 4.000 235.640 311.970 247.840 ;
        RECT 4.000 234.240 311.570 235.640 ;
        RECT 4.000 215.240 311.970 234.240 ;
        RECT 4.400 213.840 311.970 215.240 ;
        RECT 4.000 201.640 311.970 213.840 ;
        RECT 4.000 200.240 311.570 201.640 ;
        RECT 4.000 177.840 311.970 200.240 ;
        RECT 4.400 176.440 311.970 177.840 ;
        RECT 4.000 164.240 311.970 176.440 ;
        RECT 4.000 162.840 311.570 164.240 ;
        RECT 4.000 143.840 311.970 162.840 ;
        RECT 4.400 142.440 311.970 143.840 ;
        RECT 4.000 130.240 311.970 142.440 ;
        RECT 4.000 128.840 311.570 130.240 ;
        RECT 4.000 106.440 311.970 128.840 ;
        RECT 4.400 105.040 311.970 106.440 ;
        RECT 4.000 92.840 311.970 105.040 ;
        RECT 4.000 91.440 311.570 92.840 ;
        RECT 4.000 72.440 311.970 91.440 ;
        RECT 4.400 71.040 311.970 72.440 ;
        RECT 4.000 55.440 311.970 71.040 ;
        RECT 4.000 54.040 311.570 55.440 ;
        RECT 4.000 35.040 311.970 54.040 ;
        RECT 4.400 33.640 311.970 35.040 ;
        RECT 4.000 21.440 311.970 33.640 ;
        RECT 4.000 20.040 311.570 21.440 ;
        RECT 4.000 10.715 311.970 20.040 ;
      LAYER met4 ;
        RECT 81.255 11.735 174.240 311.265 ;
        RECT 176.640 11.735 177.540 311.265 ;
        RECT 179.940 11.735 272.025 311.265 ;
  END
END Guitar_Villains
END LIBRARY

